`define BR_BUS_LEN      33

`define IF2ID_pc        32
`define IF2ID_inst      32

`define IFReg_BUS_LEN   64

`define ID2EX_LEN       76
`define ID2MEM_LEN      37
`define ID2WB_LEN       39 

`define IDReg_BUS_LEN   152

`define EX2MEM_LEN      68
`define EX2WB_LEN       39

`define EXReg_BUS_LEN   107

`define MEM2WB_LEN      103

`define MEMReg_BUS_LEN  103