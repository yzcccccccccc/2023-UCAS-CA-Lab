/*************************************************
    Wrapper for AXI-SRAM-alike protocol and TLB.
    Created by yzcc, 2023.11.6
*************************************************/
module mmu_top(
    input   wire        clk,
    input   wire        reset
);


endmodule