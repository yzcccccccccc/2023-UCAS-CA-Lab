`define BR_BUS_LEN      33

`define IF2ID_pc        32
`define IF2ID_inst      32

`define ID2EX_LEN       66
`define ID2MEM_LEN      34
`define ID2WB_LEN       39 

`define EX2MEM_LEN      68
`define EX2WB_LEN       39

`define MEM2WB_LEN      103