/*****************************************************
            Control and State Reg File
    - version1.0
    - 2023.10.15, created by yzcc
******************************************************/

module csreg_file(
    input   wire        clk,
    input   wire        reset,
    input   wire        csr_re,         // enable
    input   wire [13:0] csr_num,        // addr
    output  wire [31:0] csr_rvalue,     // return value
    input   wire 
);

endmodule