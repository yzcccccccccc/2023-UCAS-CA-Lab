/************************************************************
    AXI-SRAM converter. For exp15 & exp16
*************************************************************/

module AXI_convert(
    // Input SRAM Signals

    // Output AXI signals
);

endmodule